`ifndef _csr_list_vh_
 `define _csr_list_vh_

 `define CSR_CYCLE 12'hC00
 `define CSR_TIME 12'hC01

`endif
