`ifndef _exception_vector_vh_
 `define _exception_vector_vh_
 `define VEC_RESET 32'h0
 `define VEC_ILLEGAL_INST 32'h4
 `define VEC_MISALIGNED 32'h8
`endif
