/*
 */
module core
  (
   );
endmodule // core
