`timescale 1ns / 1ps
`default_nettype none

module core_tb();
   `include "core/opcode.vh"
   reg clk_tb, resetb_tb;
   wire dm_we_tb;
   wire [31:0] im_addr_tb, dm_addr_tb, dm_di_tb;
   wire [31:0] im_do_tb, dm_do_tb;
   wire [3:0]  dm_be_tb;
   wire        dm_is_signed_tb;
   wire [11:2] im_addr_out_tb;
   wire [31:0] im_data_tb, io_data_read_tb, io_data_write_tb;
   wire [7:0]  io_addr_tb;
   wire        io_en_tb, io_we_tb;

   reg [31:0]  instruction_memory_tb [0:1023];

   reg [31:0]  io_memory_tb [0:255];

   integer     i;

   reg [32767:0] im_rom_flattened;
   always @ (*) begin
      for (i=0; i<1024; i=i+1) 
	im_rom_flattened[i*4+:32] = instruction_memory_tb[i];
   end

   reg [255:0] FD_disasm_opcode;
   always @ (*) begin : Disassembly
      case (UUT.inst_dec.opcode[6:2])
	`LOAD: FD_disasm_opcode = "LOAD    ";
	`OP_IMM: begin
	   case (UUT.inst_dec.funct3)
	     3'b000: FD_disasm_opcode = "ADDI    ";
	     3'b001: FD_disasm_opcode = "SLLI    ";
	     3'b010: FD_disasm_opcode = "SLTI    ";
	     3'b011: FD_disasm_opcode = "SLTIU   ";
	     3'b100: FD_disasm_opcode = "XORI    ";
	     3'b101: FD_disasm_opcode = UUT.inst_dec.funct7[5] 
					? "SRAI    " : "SRLI    ";
	     3'b110: FD_disasm_opcode = "ORI     ";
	     3'b111: FD_disasm_opcode = "ANDI    ";
	     default: FD_disasm_opcode = "OP-IMM  ";
	   endcase
	end
	`AUIPC: FD_disasm_opcode = "AUIPC   ";
	`STORE: FD_disasm_opcode = "STORE   ";
	`OP: begin
	   case (UUT.inst_dec.funct3)
	     3'b000: FD_disasm_opcode = UUT.inst_dec.funct7[5] ? "SUB     " : "ADD     ";
	     3'b001: FD_disasm_opcode = "SLL     ";
	     3'b010: FD_disasm_opcode = "SLT     ";
	     3'b011: FD_disasm_opcode = "SLTU    ";
	     3'b100: FD_disasm_opcode = "XOR     ";
	     3'b101: FD_disasm_opcode = UUT.inst_dec.funct7[5] ? "SRA     " : "SRL     ";
	     3'b110: FD_disasm_opcode = "OR      ";
	     3'b111: FD_disasm_opcode = "AND     ";
	     default: 	   FD_disasm_opcode = "OP?     ";
	   endcase
	end
	`LUI:  FD_disasm_opcode = "LUI     ";
	`BRANCH: FD_disasm_opcode = "BRANCH  ";
	`JALR: FD_disasm_opcode = "JALR    ";
	`JAL: FD_disasm_opcode = "JAL     ";
	`SYSTEM: FD_disasm_opcode = "SYSTEM  ";
	default: FD_disasm_opcode = "ILLEGAL ";
      endcase
   end

   always begin : CLK_GENERATOR
      #5 clk_tb = 1'b0;
      #5 clk_tb = 1'b1;
   end

   task hard_reset;
      begin
	 resetb_tb = 1'b0;
	 @(posedge clk_tb) resetb_tb = 1'b1;
      end
   endtask // hard_reset

   task load_program;
      input [2047:0] path;
      integer 	     fid, tmp;
      reg [7:0]      bytes [0:4095];
      integer 	     i,j;
      begin
	 // Initialize the instruction memory and io memory for testing
	 fid = $fopen(path, "rb");
	 tmp = $fread(bytes, fid);
	 $fclose(fid);
	 for (i=0; i<1024; i=i+1) begin
	    for (j=0; j<4; j=j+1) begin
	       instruction_memory_tb[i][8*j+:8] = bytes[i*4+j];
	    end
	 end
      end
   endtask // load_program

   task render_pipeline;
      begin
      end
   endtask

   // Test 0: NOP
   task run_test0;
      integer 	    i;
      begin
	 $display("(TT) --------------------------------------------------");
	 $display("(TT) Test 0: NOP and J Test ");
	 $display("(TT) 1. Waveform must be inspected");
	 $display("(TT) 2. Before reset, PC is at 0xFFFFFFFC.");
	 $display("(TT) 3. Reset PC is 0x0, which then jumps to 0xC.");
	 $display("(TT) 4. Then, increments at steps of 0x4.");
	 $display("(TT) 5. Then, jumps to 0xC after 0x20.");
	 $display("(TT) --------------------------------------------------");

	 load_program("tb_out/00-nop.bin");
	 hard_reset();
	 for (i=0; i<16; i=i+1) begin
	    $display("(TT) Opcode=%s, FD_PC=0x%h", FD_disasm_opcode, UUT.FD_PC);
	    @(posedge clk_tb);
	 end
      end	 
   endtask //

   // Test 1: OP-IMM
   task run_test1;
      integer 	    i;
      begin
	 $display("(TT) --------------------------------------------------");
	 $display("(TT) Test 1: OP-IMM Test ");
	 $display("(TT) 1. Waveform must be inspected");
	 $display("(TT) 2. OP-IMM's start at PC=10, depositing x1 in XB stage");
	 $display("(TT) 3. x1=1,2,3,4,5,6,1,2,1,0,1,-1,-1");
	 $display("(TT) 4. Loops to 0x0C at 0x40");
	 $display("(TT) --------------------------------------------------");

	 load_program("tb_out/01-opimm.bin");
	 hard_reset();
	 for (i=0; i<20; i=i+1) begin
	    $display("(TT) Opcode=%s, FD_PC=0x%h, x1=0x%h", 
		     FD_disasm_opcode, UUT.FD_PC, UUT.RF.data[1]);
	    @(posedge clk_tb);
	 end
      end	 
   endtask //

   // Test 2: OP-IMM
   task run_test2;
      integer 	    i;
      begin
	 $display("(TT) --------------------------------------------------");
	 $display("(TT) Test 2: OP Test ");
	 $display("(TT) 1. Waveform must be inspected");
	 $display("(TT) 2. OP's start at PC=14. x1 has 2 clock delay");
	 $display("(TT) 3. x1=4,3,1,0,1,0,1,2,4,2,-2,-1,1,0,1");
	 $display("(TT) 4. Loops to 0x0C at 50");
	 $display("(TT) --------------------------------------------------");

	 load_program("tb_out/02-op.bin");
	 hard_reset();
	 for (i=0; i<24; i=i+1) begin
	    $display("(TT) Opcode=%s, FD_PC=0x%h, x1=0x%h", 
		     FD_disasm_opcode, UUT.FD_PC, UUT.RF.data[1]);
	    @(posedge clk_tb);
	 end
      end	 
   endtask //
   
   assign im_data_tb = instruction_memory_tb[im_addr_out_tb[11:2]];
   assign io_data_read_tb = io_memory_tb[io_addr_tb[7:2]];
   
   mmu MMU0(.clk(clk_tb), .resetb(resetb_tb), .dm_we(dm_we_tb), 
	   .im_addr(im_addr_tb), .im_do(im_do_tb),
	   .dm_addr(dm_addr_tb), .dm_di(dm_di_tb),
	   .dm_do(dm_do_tb), .dm_be(dm_be_tb),
	   .is_signed(dm_is_signed_tb),
	   .im_addr_out(im_addr_out_tb), .im_data(im_data_tb),
	   .io_addr(io_addr_tb), .io_en(io_en_tb), .io_we(io_we_tb),
	   .io_data_read(io_data_read_tb), .io_data_write(io_data_write_tb)
	   );

   core UUT
     (
      .clk(clk_tb), .resetb(resetb_tb),
      .dm_we(dm_we_tb), .im_addr(im_addr_tb),
      .im_do(im_do_tb), .dm_addr(dm_addr_tb),
      .dm_di(dm_di_tb), .dm_do(dm_do_tb),
      .dm_be(dm_be_tb), .dm_is_signed(dm_is_signed_tb)
      );

   // Run the tests
   initial
     begin : RUN_ALL_TESTS
	$dumpfile("tb_log/core_tb.vcd");
	$dumpvars(0,core_tb);
	for (i = 0; i < 256; i = i + 1) begin
	   io_memory_tb[i] = 4096 + i;
	end

	@(posedge clk_tb);

	run_test0();
	run_test1();
	run_test2();

	$finish;
	
     end


endmodule 

