`ifndef _exception_vector_vh_
 `define _exception_vector_vh_
 `define VEC_RESET 32'h0
 `define VEC_DEFAULT 32'h4
`endif
