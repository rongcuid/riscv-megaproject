`ifndef _aluop_vh_
 `define _aluop_vh_

 `define ALUOP1_UNKN 32'bX
 `define ALUOP1_RS1 0
 `define ALUOP1_PC 1

 `define ALUOP2_UNKN 32'bX
 `define ALUOP2_RS2 0
 `define ALUOP2_IMM 1

 `define ALU_UNKN 32'bX
 `define ALU_ADD 0
 `define ALU_SLT 1
 `define ALU_AND 2
 `define ALU_OR 3
 `define ALU_XOR 4
 `define ALU_SLL 5
 `define ALU_SRL 6
 `define ALU_SRA 7
 `define ALU_SUB 8

`endif
